`timescale 1ns / 1ps

module instr_fetcher(
	input [31:0] pc,
	input clk,
	output [31:0] instr
   );
	
	instructions 


endmodule
